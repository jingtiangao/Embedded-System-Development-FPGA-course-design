DFF1.VHD,FADDER.VHD)
FBRAC.VHD
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY FBRAC IS
  PORT( aT:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		bT:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		sT:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		CINTOP:IN STD_LOGIC;
		CLKTOP :IN STD_LOGIC;
		COUTTOP : OUT STD_LOGIC);
END ENTITY FBRAC;
ARCHITECTURE ONE OF FBRAC IS
COMPONENT DFF1
 PORT (D:IN STD_LOGIC;
	   CLK:IN STD_LOGIC;
	   Q:OUT STD_LOGIC);
END COMPONENT DFF1;

COMPONENT RFF1
 PORT(CLK :IN STD_LOGIC;
	  R :  IN STD_LOGIC_VECTOR(3 DOWNTO 0);	
	  Q :  OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END COMPONENT RFF1;
COMPONENT bit4_f_adder
PORT(aa:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	 bb:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	 cin:IN STD_LOGIC;
	 cout:OUT STD_LOGIC;
	 ss:OUT STD_LOGIC_VECTOR(3 DOWNTO 0));

END COMPONENT bit4_f_adder;
SIGNAL E,F,G: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL D1 :STD_LOGIC;
BEGIN
U1: RFF1 PORT MAP(R=>aT,Q=>E,CLK=>CLKTOP);
U2: RFF1 PORT MAP(R=>bT,Q=>F,CLK=>CLKTOP);
U3: bit4_f_adder PORT MAP(aa=>E,bb=>F,cin=>CINTOP,cout=>D1,ss=>G);
U4: RFF1 PORT MAP(R=>G,Q=>sT,CLK=>CLKTOP);
U5: DFF1 PORT MAP(D=>D1,Q=>COUTTOP,CLK=>CLKTOP);
END ARCHITECTURE ONE;
DFF1.VHD
LIBRARY IEEE ;
USE IEEE.STD_LOGIC_1164.ALL ;
ENTITY DFF1 IS
  PORT (CLK : IN STD_LOGIC ;
		  D : IN STD_LOGIC ;
		  Q : OUT STD_LOGIC );
 END ;
ARCHITECTURE bhv OF DFF1 IS
  SIGNAL Q1 : STD_LOGIC ;
  BEGIN 
   PROCESS (CLK)
	BEGIN
	 IF CLK'EVENT AND CLK = '1'
		THEN Q1 <= D ;
	 END IF ;
	    Q <= Q1;
   END PROCESS ;
END bhv ;
RFF1.VHD
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY RFF1 IS
 PORT(CLK :IN STD_LOGIC;
	  R :  IN STD_LOGIC_VECTOR(3 DOWNTO 0);	
	  Q :  OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END ENTITY RFF1;
ARCHITECTURE rhv OF RFF1 IS
	SIGNAL A: STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN
	  PROCESS(CLK)
	  BEGIN
	   IF CLK'EVENT AND CLK ='1'
		  THEN  A<= R;
	   END IF;
		Q<= A;

	  END PROCESS ;
END rhv;
bit4_f_adder.VHD
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY bit4_f_adder IS
  PORT(aa : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
       bb : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
       cin: IN STD_LOGIC;
       cout: OUT STD_LOGIC;
       ss : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END ENTITY bit4_f_adder;

ARCHITECTURE one OF bit4_f_adder IS
  COMPONENT f_adder
    PORT (a, b, c: IN STD_LOGIC;
           CO, SO: OUT STD_LOGIC);
    END COMPONENT;
  SIGNAL C1, C2, C3: STD_LOGIC;
  BEGIN
    U1 : f_adder PORT MAP(c=>cin, a=>aa(0), b=>bb(0), SO=>ss(0), CO=>C1 );
    U2 : f_adder PORT MAP(c=>C1, a=>aa(1), b=>bb(1), SO=>ss(1), CO=>C2 );
    U3 : f_adder PORT MAP(c=>C2, a=>aa(2), b=>bb(2), SO=>ss(2), CO=>C3 );
    U4 : f_adder PORT MAP(c=>C3, a=>aa(3), b=>bb(3), SO=>ss(3), CO=>cout );
END ARCHITECTURE one;
f_adder.VHD
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY f_adder IS 
  PORT (a, b, c: IN STD_LOGIC;
           CO, SO: OUT STD_LOGIC);
END ENTITY f_adder;

ARCHITECTURE one OF f_adder IS
   SIGNAL abc : STD_LOGIC_VECTOR(2 DOWNTO 0);
   SIGNAL CSO : STD_LOGIC_VECTOR(1 DOWNTO 0);
   BEGIN 
      abc <= a&b&c;
   PROCESS(abc)
   BEGIN 
      CASE abc IS
      WHEN "000" => CSO <= "00";
      WHEN "010" => CSO <= "01";
      WHEN "100" => CSO <= "01";
      WHEN "110" => CSO <= "10";
      WHEN "001" => CSO <= "01";
      WHEN "011" => CSO <= "10";
      WHEN "101" => CSO <= "10";
      WHEN "111" => CSO <= "11";
      WHEN OTHERS => NULL;
      END CASE;
   
   END PROCESS;
   CO<=CSO(1);SO<=CSO(0);
END ARCHITECTURE one;	
